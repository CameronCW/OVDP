// OVDP.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module OVDP (
		input  wire       clk_clk,                              //                            clk.clk
		output wire       i2s_tx_bclk_export,                   //                    i2s_tx_bclk.export
		output wire       i2s_tx_lrclk_export,                  //                   i2s_tx_lrclk.export
		output wire       i2s_tx_sdata_export,                  //                   i2s_tx_sdata.export
		output wire [7:0] pid_focus_pwm_out_export,             //              pid_focus_pwm_out.export
		input  wire       preprocess_block_lsync_export,        //         preprocess_block_lsync.export
		input  wire       preprocess_block_rsync_export,        //         preprocess_block_rsync.export
		input  wire       preprocess_block_sig_export,          //           preprocess_block_sig.export
		input  wire       reset_reset_n,                        //                          reset.reset_n
		input  wire       spislave_avalon_streaming_sink_valid, // spislave_avalon_streaming_sink.valid
		input  wire [7:0] spislave_avalon_streaming_sink_data,  //                               .data
		output wire       spislave_avalon_streaming_sink_ready, //                               .ready
		input  wire       spislave_export_mosi,                 //                spislave_export.mosi
		input  wire       spislave_export_nss,                  //                               .nss
		inout  wire       spislave_export_miso,                 //                               .miso
		input  wire       spislave_export_sclk                  //                               .sclk
	);

	wire         pll_0_outclk0_clk;                         // pll_0:outclk_0 -> [channel_processor_top_0:clk_slow, pid_focus_0:clk_slow]
	wire         preprocess_block_0_dir_export;             // preProcess_block_0:dir -> sig_extract_0:dir
	wire         preprocess_block_0_dir_cp_export;          // preProcess_block_0:dir_cp -> channel_processor_top_0:dir
	wire  [15:0] spi_command_decoder_0_focus_signal_export; // spi_command_decoder_0:focus_signal -> pid_focus_0:focus_signal
	wire  [15:0] spi_command_decoder_0_kd_export;           // spi_command_decoder_0:kd -> pid_focus_0:kd
	wire  [15:0] spi_command_decoder_0_ki_export;           // spi_command_decoder_0:ki -> pid_focus_0:ki
	wire  [15:0] spi_command_decoder_0_kp_export;           // spi_command_decoder_0:kp -> pid_focus_0:kp
	wire         spi_command_decoder_0_mute_export;         // spi_command_decoder_0:mute -> output_conversion_0:mute
	wire  [15:0] output_conversion_0_out_l_export;          // output_conversion_0:out_L -> i2s_tx_0:sample_L
	wire  [15:0] output_conversion_0_out_r_export;          // output_conversion_0:out_R -> i2s_tx_0:sample_R
	wire  [15:0] channel_processor_top_0_sample_l_export;   // channel_processor_top_0:sample_L -> output_conversion_0:sample_L
	wire  [15:0] channel_processor_top_0_sample_r_export;   // channel_processor_top_0:sample_R -> output_conversion_0:sample_R
	wire         sig_extract_0_sample_pair_valid_export;    // sig_extract_0:sample_pair_valid -> channel_processor_top_0:sample_valid
	wire         preprocess_block_0_sig_fall_l_export;      // preProcess_block_0:sig_fall_L -> sig_extract_0:sig_fall_L
	wire         preprocess_block_0_sig_fall_r_export;      // preProcess_block_0:sig_fall_R -> sig_extract_0:sig_fall_R
	wire         preprocess_block_0_sig_rise_l_export;      // preProcess_block_0:sig_rise_L -> sig_extract_0:sig_rise_L
	wire         preprocess_block_0_sig_rise_r_export;      // preProcess_block_0:sig_rise_R -> sig_extract_0:sig_rise_R
	wire  [31:0] sig_extract_0_left_sample_time_export;     // sig_extract_0:left_sample_time -> channel_processor_top_0:sig_time_L
	wire  [31:0] preprocess_block_0_sig_time_l_export;      // preProcess_block_0:sig_time_L -> sig_extract_0:sig_time_L
	wire  [31:0] sig_extract_0_right_sample_time_export;    // sig_extract_0:right_sample_time -> channel_processor_top_0:sig_time_R
	wire  [31:0] preprocess_block_0_sig_time_r_export;      // preProcess_block_0:sig_time_R -> sig_extract_0:sig_time_R
	wire  [31:0] preprocess_block_0_split_sync_time_export; // preProcess_block_0:split_sync_time -> sig_extract_0:split_sync_time
	wire         preprocess_block_0_sync_start_export;      // preProcess_block_0:sync_start -> channel_processor_top_0:sync_start
	wire  [31:0] preprocess_block_0_t_ltr_export;           // preProcess_block_0:t_ltr -> channel_processor_top_0:t_ltr
	wire  [31:0] preprocess_block_0_t_rtl_export;           // preProcess_block_0:t_rtl -> channel_processor_top_0:t_rtl
	wire  [15:0] spi_command_decoder_0_threshold_export;    // spi_command_decoder_0:threshold -> pid_focus_0:threshold
	wire         channel_processor_top_0_valid_l_export;    // channel_processor_top_0:valid_L -> output_conversion_0:valid_L
	wire         channel_processor_top_0_valid_r_export;    // channel_processor_top_0:valid_R -> output_conversion_0:valid_R
	wire         output_conversion_0_valid_out_export;      // output_conversion_0:valid_out -> i2s_tx_0:valid_in
	wire   [7:0] spi_command_decoder_0_volume_export;       // spi_command_decoder_0:volume -> output_conversion_0:volume
	wire         spislave_0_avalon_streaming_source_valid;  // spislave_0:stsourcevalid -> avalon_st_adapter:in_0_valid
	wire   [7:0] spislave_0_avalon_streaming_source_data;   // spislave_0:stsourcedata -> avalon_st_adapter:in_0_data
	wire         spislave_0_avalon_streaming_source_ready;  // avalon_st_adapter:in_0_ready -> spislave_0:stsourceready
	wire         avalon_st_adapter_out_0_valid;             // avalon_st_adapter:out_0_valid -> spi_command_decoder_0:stream_valid
	wire   [7:0] avalon_st_adapter_out_0_data;              // avalon_st_adapter:out_0_data -> spi_command_decoder_0:stream_data
	wire         rst_controller_reset_out_reset;            // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, channel_processor_top_0:reset_n, i2s_tx_0:reset_n, output_conversion_0:reset_n, pid_focus_0:reset_n, preProcess_block_0:reset_n, sig_extract_0:reset_n, spi_command_decoder_0:reset_n, spislave_0:nreset]

	channel_processor_top channel_processor_top_0 (
		.clk          (clk_clk),                                 //        clock.clk
		.reset_n      (~rst_controller_reset_out_reset),         //        reset.reset_n
		.sample_L     (channel_processor_top_0_sample_l_export), //     sample_L.export
		.sample_R     (channel_processor_top_0_sample_r_export), //     sample_R.export
		.sample_valid (sig_extract_0_sample_pair_valid_export),  // sample_valid.export
		.sig_time_L   (sig_extract_0_left_sample_time_export),   //   sig_time_L.export
		.sig_time_R   (sig_extract_0_right_sample_time_export),  //   sig_time_R.export
		.sync_start   (preprocess_block_0_sync_start_export),    //   sync_start.export
		.t_ltr        (preprocess_block_0_t_ltr_export),         //        t_ltr.export
		.t_rtl        (preprocess_block_0_t_rtl_export),         //        t_rtl.export
		.valid_L      (channel_processor_top_0_valid_l_export),  //      valid_L.export
		.valid_R      (channel_processor_top_0_valid_r_export),  //      valid_R.export
		.dir          (preprocess_block_0_dir_cp_export),        //          dir.export
		.clk_slow     (pll_0_outclk0_clk)                        //   clock_slow.clk
	);

	i2s_transmitter i2s_tx_0 (
		.clk      (clk_clk),                              //    clock.clk
		.reset_n  (~rst_controller_reset_out_reset),      //    reset.reset_n
		.valid_in (output_conversion_0_valid_out_export), // valid_in.export
		.sdata    (i2s_tx_sdata_export),                  //    sdata.export
		.sample_L (output_conversion_0_out_l_export),     // sample_L.export
		.sample_R (output_conversion_0_out_r_export),     // sample_R.export
		.lrclk    (i2s_tx_lrclk_export),                  //    lrclk.export
		.bclk     (i2s_tx_bclk_export)                    //     bclk.export
	);

	output_conversion output_conversion_0 (
		.clk       (clk_clk),                                 //     clock.clk
		.reset_n   (~rst_controller_reset_out_reset),         //     reset.reset_n
		.mute      (spi_command_decoder_0_mute_export),       //      mute.export
		.out_R     (output_conversion_0_out_r_export),        //     out_R.export
		.sample_L  (channel_processor_top_0_sample_l_export), //  sample_L.export
		.sample_R  (channel_processor_top_0_sample_r_export), //  sample_R.export
		.valid_L   (channel_processor_top_0_valid_l_export),  //   valid_L.export
		.valid_R   (channel_processor_top_0_valid_r_export),  //   valid_R.export
		.valid_out (output_conversion_0_valid_out_export),    // valid_out.export
		.volume    (spi_command_decoder_0_volume_export),     //    volume.export
		.out_L     (output_conversion_0_out_l_export)         //     out_L.export
	);

	pid_focus_controller pid_focus_0 (
		.clk          (clk_clk),                                   //        clock.clk
		.reset_n      (~rst_controller_reset_out_reset),           //        reset.reset_n
		.focus_signal (spi_command_decoder_0_focus_signal_export), // focus_signal.export
		.kp           (spi_command_decoder_0_kp_export),           //           kp.export
		.ki           (spi_command_decoder_0_ki_export),           //           ki.export
		.kd           (spi_command_decoder_0_kd_export),           //           kd.export
		.pwm_out      (pid_focus_pwm_out_export),                  //      pwm_out.export
		.threshold    (spi_command_decoder_0_threshold_export),    //    threshold.export
		.clk_slow     (pll_0_outclk0_clk)                          //   clock_slow.clk
	);

	OVDP_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

	preprocess_block preprocess_block_0 (
		.clk             (clk_clk),                                   //           clock.clk
		.reset_n         (~rst_controller_reset_out_reset),           //           reset.reset_n
		.dir             (preprocess_block_0_dir_export),             //             dir.export
		.lsync           (preprocess_block_lsync_export),             //           lsync.export
		.rsync           (preprocess_block_rsync_export),             //           rsync.export
		.sig             (preprocess_block_sig_export),               //             sig.export
		.sig_fall_L      (preprocess_block_0_sig_fall_l_export),      //      sig_fall_L.export
		.sig_fall_R      (preprocess_block_0_sig_fall_r_export),      //      sig_fall_R.export
		.sig_rise_L      (preprocess_block_0_sig_rise_l_export),      //      sig_rise_L.export
		.sig_rise_R      (preprocess_block_0_sig_rise_r_export),      //      sig_rise_R.export
		.sig_time_L      (preprocess_block_0_sig_time_l_export),      //      sig_time_L.export
		.split_sync_time (preprocess_block_0_split_sync_time_export), // split_sync_time.export
		.sync_start      (preprocess_block_0_sync_start_export),      //      sync_start.export
		.t_ltr           (preprocess_block_0_t_ltr_export),           //           t_ltr.export
		.t_rtl           (preprocess_block_0_t_rtl_export),           //           t_rtl.export
		.sig_time_R      (preprocess_block_0_sig_time_r_export),      //      sig_time_R.export
		.dir_cp          (preprocess_block_0_dir_cp_export)           //          dir_cp.export
	);

	sig_extract sig_extract_0 (
		.clk               (clk_clk),                                   //             clock.clk
		.reset_n           (~rst_controller_reset_out_reset),           //             reset.reset_n
		.split_sync_time   (preprocess_block_0_split_sync_time_export), //   split_sync_time.export
		.dir               (preprocess_block_0_dir_export),             //               dir.export
		.left_sample_time  (sig_extract_0_left_sample_time_export),     //  left_sample_time.export
		.right_sample_time (sig_extract_0_right_sample_time_export),    // right_sample_time.export
		.sample_pair_valid (sig_extract_0_sample_pair_valid_export),    // sample_pair_valid.export
		.sig_fall_L        (preprocess_block_0_sig_fall_l_export),      //        sig_fall_L.export
		.sig_fall_R        (preprocess_block_0_sig_fall_r_export),      //        sig_fall_R.export
		.sig_rise_L        (preprocess_block_0_sig_rise_l_export),      //        sig_rise_L.export
		.sig_rise_R        (preprocess_block_0_sig_rise_r_export),      //        sig_rise_R.export
		.sig_time_L        (preprocess_block_0_sig_time_l_export),      //        sig_time_L.export
		.sig_time_R        (preprocess_block_0_sig_time_r_export)       //        sig_time_R.export
	);

	spi_command_decoder spi_command_decoder_0 (
		.clk          (clk_clk),                                   //                 clock.clk
		.reset_n      (~rst_controller_reset_out_reset),           //                 reset.reset_n
		.stream_data  (avalon_st_adapter_out_0_data),              // avalon_streaming_sink.data
		.stream_valid (avalon_st_adapter_out_0_valid),             //                      .valid
		.ki           (spi_command_decoder_0_ki_export),           //                    ki.export
		.kp           (spi_command_decoder_0_kp_export),           //                    kp.export
		.kd           (spi_command_decoder_0_kd_export),           //                    kd.export
		.mute         (spi_command_decoder_0_mute_export),         //                  mute.export
		.focus_signal (spi_command_decoder_0_focus_signal_export), //          focus_signal.export
		.threshold    (spi_command_decoder_0_threshold_export),    //             threshold.export
		.volume       (spi_command_decoder_0_volume_export)        //                volume.export
	);

	SPIPhy #(
		.SYNC_DEPTH (3)
	) spislave_0 (
		.sysclk        (clk_clk),                                  //              clock_sink.clk
		.nreset        (~rst_controller_reset_out_reset),          //        clock_sink_reset.reset_n
		.mosi          (spislave_export_mosi),                     //                export_0.export
		.nss           (spislave_export_nss),                      //                        .export
		.miso          (spislave_export_miso),                     //                        .export
		.sclk          (spislave_export_sclk),                     //                        .export
		.stsourceready (spislave_0_avalon_streaming_source_ready), // avalon_streaming_source.ready
		.stsourcevalid (spislave_0_avalon_streaming_source_valid), //                        .valid
		.stsourcedata  (spislave_0_avalon_streaming_source_data),  //                        .data
		.stsinkvalid   (spislave_avalon_streaming_sink_valid),     //   avalon_streaming_sink.valid
		.stsinkdata    (spislave_avalon_streaming_sink_data),      //                        .data
		.stsinkready   (spislave_avalon_streaming_sink_ready)      //                        .ready
	);

	OVDP_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (0),
		.inDataWidth     (8),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (0),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk   (clk_clk),                                  // in_clk_0.clk
		.in_rst_0_reset (rst_controller_reset_out_reset),           // in_rst_0.reset
		.in_0_data      (spislave_0_avalon_streaming_source_data),  //     in_0.data
		.in_0_valid     (spislave_0_avalon_streaming_source_valid), //         .valid
		.in_0_ready     (spislave_0_avalon_streaming_source_ready), //         .ready
		.out_0_data     (avalon_st_adapter_out_0_data),             //    out_0.data
		.out_0_valid    (avalon_st_adapter_out_0_valid)             //         .valid
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
